Version 4
SHEET 1 896 680
WIRE -48 -16 -64 -16
WIRE 48 -16 32 -16
WIRE 112 -16 48 -16
WIRE 208 -16 192 -16
WIRE 112 64 112 48
WIRE 48 80 48 -16
WIRE 80 80 48 80
WIRE 208 96 208 -16
WIRE 208 96 144 96
WIRE -400 112 -400 80
WIRE -272 112 -272 80
WIRE 80 112 -16 112
WIRE -16 144 -16 112
WIRE 112 144 112 128
WIRE -400 240 -400 192
WIRE -272 240 -272 192
WIRE -16 256 -16 224
FLAG -272 240 0
FLAG 112 48 +V
FLAG -272 80 +V
FLAG 112 144 -V
FLAG -400 240 0
FLAG -400 80 -V
FLAG -16 256 0
FLAG -64 -16 0
SYMBOL voltage -272 96 R0
SYMATTR InstName V1
SYMATTR Value 2.5
SYMBOL voltage -400 96 R0
SYMATTR InstName V2
SYMATTR Value -2.5
SYMBOL voltage -16 128 R0
SYMATTR InstName V3
SYMATTR Value SINE(0 1 1K)
SYMBOL res 208 -32 R90
WINDOW 0 0 56 VBottom 2
WINDOW 3 32 56 VTop 2
SYMATTR InstName R1
SYMATTR Value 10K
SYMBOL res 48 -32 R90
WINDOW 0 0 56 VBottom 2
WINDOW 3 32 56 VTop 2
SYMATTR InstName R2
SYMATTR Value 10K
SYMBOL LTC2055 112 96 R0
SYMATTR InstName U1
TEXT -192 296 Left 2 !.tran 3m
